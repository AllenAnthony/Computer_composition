// Verilog test fixture created from schematic E:\ISE\work\multy_CPU\top_for_multy_CPU.sch - Sun Jun 12 21:20:44 2016

`timescale 1ns / 1ps

module top_for_multy_CPU_top_for_multy_CPU_sch_tb();

// Inputs
   reg clk;
   reg [4:0] SW;

// Output

// Bidirs

// Instantiate the UUT
   top_for_multy_CPU UUT (
		.clk(clk), 
		.SW(SW)
   );
// Initialize Inputs
   
   
endmodule
